module example_crg_inst(
input clk,
input rst_n);
wire    clk_phy_en;
wire    clk_phy;
wire    rst_clk_phy;
wire    clk1_sel;
wire    clk1_en;
wire    clk1;
wire    rst_clk1;
wire    clk2_en;
wire    clk2;
wire    rst_clk2;
wire    clk3_en;
wire    clk3;
wire    rst_clk3;
example_crg u_crg(
    .clk_phy_en                         (clk_phy_en),
   .clk_phy                             (clk_phy),
   .rst_clk_phy                         (rst_clk_phy),
    .clk1_sel                           (clk1_sel),
    .clk1_en                            (clk1_en),
   .clk1                                (clk1),
   .rst_clk1                            (rst_clk1),
    .clk2_en                            (clk2_en),
   .clk2                                (clk2),
   .rst_clk2                            (rst_clk2),
    .clk3_en                            (clk3_en),
   .clk3                                (clk3),
   .rst_clk3                            (rst_clk3),
   .clk_src                             (ap_clk),
   .rst_n_sys                           (ap_rst_n));
endmodule