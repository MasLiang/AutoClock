module module_1_crg_inst(
input clk,
input rst_n);
wire    clk1_sel;
wire    clk1_en;
wire    clk1;
wire    rst_clk1;
wire    clk3_en;
wire    clk3;
wire    rst_clk3;
module_1_crg u_crg(
    .clk1_sel                           (clk1_sel),
    .clk1_en                            (clk1_en),
   .clk1                                (clk1),
   .rst_clk1                            (rst_clk1),
    .clk3_en                            (clk3_en),
   .clk3                                (clk3),
   .rst_clk3                            (rst_clk3),
   .clk_src                             (ap_clk),
   .rst_n_sys                           (ap_rst_n));
endmodule